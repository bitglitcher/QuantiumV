module regfile();
  
  
  
endmodule
