module d_cache();
  
  
  
endmodule
