module fetch_stage();



emdmodule
