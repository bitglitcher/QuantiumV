// SPDX-License-Identifier: MIT

/* This file contains the defaults for Wishbone. */

/* ------------------------------------------------------------------------- */


// TODO


/* ------------------------------------------------------------------------- */


/* End of file. */
