module soc();
  
  
  
endmodule
