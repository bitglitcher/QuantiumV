module alu();
  
  
  
endmodule
