module core
  (
    input clk,
    input rst
  );
  
  
  
  
  
endmodule
