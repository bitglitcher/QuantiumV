module i_cache();



endmodule
