// SPDX-License-Identifier: MIT

/* This file contains the defaults for AXI. */

/* ------------------------------------------------------------------------- */


// TODO


/* ------------------------------------------------------------------------- */


/* End of file. */
